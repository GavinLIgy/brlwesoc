module tb_user_ram()



endmodule